-- global package

library IEEE;
use IEEE.std_logic_1164.all;

package my_pkg is

	type sixteenbyeight is array (15 downto 0) of std_logic_vector(7 downto 0);

	
end my_pkg;